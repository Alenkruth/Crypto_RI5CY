`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Engineer:     Alenkruth                                                    //
// Project:      RISC-V crypto Extension                                      //
//                               //
////////////////////////////////////////////////////////////////////////////////


module riscv_c_test(

    );
endmodule
